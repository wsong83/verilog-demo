
// 多功能计算器
module (
  input [3:0] a, b,
  input [2:0] s,
  output [4:0] y);

// 下面是计算机的内部实现代码





endmodule


